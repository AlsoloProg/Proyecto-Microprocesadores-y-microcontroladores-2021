`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/15/2021 11:11:39 PM
// Design Name: 
// Module Name: MemInstru
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module MemInstru (Direccion, B1, B2, B3, B4); // Memoria de instrucciones
    
    input [6:0] Direccion; // entra PC

    reg [7:0] ROMINSTRU [127:0]; // se inicializa la memoria con 128 espacios de 8 bits c/u
    output reg [7:0] B1; // salen los bits m�s significativos de la instrucci�n
    output reg [7:0] B2; // salen los siguientes cuatro bits de la instrucci�n
    output reg [7:0] B3; // salen los siguientes cuatro bits de la instrucci�n
    output reg [7:0] B4; // salen los bits menos significativos de la instrucci�n
   
    initial begin
        $readmemb("WhileBin.txt", ROMINSTRU); // se carga la memoria con el c�digo whilebin
    end
        
    always @(*) // se asignan las salidas de acuerdo a la direcci�n en memoria
        begin
            B1 <= ROMINSTRU[Direccion]; 
            B2 <= ROMINSTRU[Direccion+2'd1];
            B3 <= ROMINSTRU[Direccion+2'd2];
            B4 <= ROMINSTRU[Direccion+2'd3];
        end
endmodule
